library verilog;
use verilog.vl_types.all;
entity tb_mru is
end tb_mru;
